module simple_axi_master (
    input  clk,
    input  rst,
    output out
);

endmodule
